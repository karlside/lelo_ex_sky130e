magic
tech sky130A
magscale 1 2
timestamp 1769092861
<< locali >>
rect 161 1956 565 2049
rect -96 -200 96 152
rect -203 -202 400 -200
rect -203 -382 294 -202
rect 1056 -207 1248 156
rect 474 -382 1407 -207
rect -203 -399 1407 -382
rect -203 -400 400 -399
<< viali >>
rect 294 -382 474 -202
<< metal1 >>
rect 160 137 224 3900
rect 288 -202 480 3860
rect 672 3658 1143 3850
rect 951 3078 1143 3658
rect 707 2886 1143 3078
rect 951 1467 1143 2886
rect 702 1275 1143 1467
rect 951 379 1143 1275
rect 697 187 1143 379
rect 672 40 864 120
rect 288 -382 294 -202
rect 474 -382 480 -202
rect 288 -394 480 -382
use JNWATR_NCH_4C5F0  xo0<0> ../JNW_ATR_SKY130A
timestamp 1740610800
transform 1 0 0 0 1 0
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo0<1>
timestamp 1740610800
transform 1 0 0 0 1 800
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo1
timestamp 1740610800
transform 1 0 0 0 1 1600
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo2<0>
timestamp 1740610800
transform 1 0 0 0 1 2400
box -184 -128 1336 928
use JNWATR_NCH_4C5F0  xo2<1>
timestamp 1740610800
transform 1 0 0 0 1 3200
box -184 -128 1336 928
<< labels >>
flabel metal1 s 288 600 480 680 0 FreeSans 400 0 0 0 VSS
port 1 nsew ground bidirectional
flabel metal1 s 160 360 224 440 0 FreeSans 400 0 0 0 IBPS_5U
port 2 nsew signal bidirectional
flabel metal1 s 672 40 864 120 0 FreeSans 400 0 0 0 IBNS_20U
port 3 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1152 4000
<< end >>
